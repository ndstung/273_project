package project ; //user's package

    import uvm_pkg::*; //necessary to include this package in user's package
    
    
    `include "sequence_item.sv"
    `include "sequence.sv"
    `include "sequencer.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "reference.sv"
    `include "agent.sv"
    `include "scoreboard.sv"
    `include "environment.sv"
    `include "test.sv"
    
    endpackage : project